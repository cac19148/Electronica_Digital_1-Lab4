module testbench();

  reg p1_1, p2_1, p3_1, p1_2, p2_2, p3_2, p1_3, p2_3, p3_3, p1_4, p2_4, p3_4,   p4_1, p5_1, p6_1, p7_1, p4_2, p5_2, p6_2, p7_2, p4_3, p5_3, p6_3, p7_3, p4_4, p5_4, p6_4, p7_4;
  wire led1_1, led1_2, led1_3, led1_4, led2_1, led2_2, led2_3, led2_4;

  gateLevel_1   G1(p1_1, p2_1, p3_1, led1_1);
  gateLevel_2   G2(p1_2, p2_2, p3_2, led1_2);
  gateLevel_3   G3(p1_3, p2_3, p3_3, led1_3);
  gateLevel_4   G4(p1_4, p2_4, p3_4, led1_4);
  
  operadores_1 OP1(p4_1, p5_1, p6_1, p7_1, led2_1);
  operadores_2 OP2(p4_2, p5_2, p6_2, p7_2, led2_2);
  operadores_3 OP3(p4_3, p5_3, p6_3, p7_3, led2_3);
  operadores_4 OP4(p4_4, p5_4, p6_4, p7_4, led2_4);

  initial begin
	$display("");
	$display("EJERCICIO 1: TABLA 1");
    $display("A B C | Y");
    $display("------|--");
    $monitor("%b %b %b | %b", p1_1, p2_1, p3_1, led1_1);
       p1_1 = 0; p2_1 = 0; p3_1 = 0;
    #1 p1_1 = 0; p2_1 = 0; p3_1 = 1;
    #1 p1_1 = 0; p2_1 = 1; p3_1 = 0;
    #1 p1_1 = 0; p2_1 = 1; p3_1 = 1;
    #1 p1_1 = 1; p2_1 = 0; p3_1 = 0;
    #1 p1_1 = 1; p2_1 = 0; p3_1 = 1;
    #1 p1_1 = 1; p2_1 = 1; p3_1 = 0;
    #1 p1_1 = 1; p2_1 = 1; p3_1 = 1;
	#1 $display("");
  end
  
  initial begin
    #10
	$display("EJERCICIO 1: TABLA 2");
    $display("A B C | Y");
    $display("------|--");
    $monitor("%b %b %b | %b", p1_2, p2_2, p3_2, led1_2);
       p1_2 = 0; p2_2 = 0; p3_2 = 0;
    #1 p1_2 = 0; p2_2 = 0; p3_2 = 1;
    #1 p1_2 = 0; p2_2 = 1; p3_2 = 0;
    #1 p1_2 = 0; p2_2 = 1; p3_2 = 1;
    #1 p1_2 = 1; p2_2 = 0; p3_2 = 0;
    #1 p1_2 = 1; p2_2 = 0; p3_2 = 1;
    #1 p1_2 = 1; p2_2 = 1; p3_2 = 0;
    #1 p1_2 = 1; p2_2 = 1; p3_2 = 1;
	#1 $display("");
  end
  
  initial begin
    #20
	$display("EJERCICIO 2: TABLA 2");
    $display("A B C | Y");
    $display("------|--");
    $monitor("%b %b %b | %b", p1_3, p2_3, p3_3, led1_3);
       p1_3 = 0; p2_3 = 0; p3_3 = 0;
    #1 p1_3 = 0; p2_3 = 0; p3_3 = 1;
    #1 p1_3 = 0; p2_3 = 1; p3_3 = 0;
    #1 p1_3 = 0; p2_3 = 1; p3_3 = 1;
    #1 p1_3 = 1; p2_3 = 0; p3_3 = 0;
    #1 p1_3 = 1; p2_3 = 0; p3_3 = 1;
    #1 p1_3 = 1; p2_3 = 1; p3_3 = 0;
    #1 p1_3 = 1; p2_3 = 1; p3_3 = 1;
	#1 $display("");
  end
  
  initial begin
    #30
	$display("EJERCICIO 2: TABLA 4");
    $display("A B C | Y");
    $display("------|--");
    $monitor("%b %b %b | %b", p1_4, p2_4, p3_4, led1_4);
       p1_4 = 0; p2_4 = 0; p3_4 = 0;
    #1 p1_4 = 0; p2_4 = 0; p3_4 = 1;
    #1 p1_4 = 0; p2_4 = 1; p3_4 = 0;
    #1 p1_4 = 0; p2_4 = 1; p3_4 = 1;
    #1 p1_4 = 1; p2_4 = 0; p3_4 = 0;
    #1 p1_4 = 1; p2_4 = 0; p3_4 = 1;
    #1 p1_4 = 1; p2_4 = 1; p3_4 = 0;
    #1 p1_4 = 1; p2_4 = 1; p3_4 = 1;
	#1 $display("");
	#1 $display("-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-");
  end
  
  initial begin
    #40
	$display("EJERCICIO 1: TABLA 3");
    $display("A B C D | Y");
    $display("--------|--");
    $monitor("%b %b %b %b | %b", p4_1, p5_1, p6_1, p7_1, led2_1);
       p4_1 = 0; p5_1 = 0; p6_1 = 0; p7_1 = 0;
    #1 p4_1 = 0; p5_1 = 0; p6_1 = 0; p7_1 = 1;
    #1 p4_1 = 0; p5_1 = 0; p6_1 = 1; p7_1 = 0;
    #1 p4_1 = 0; p5_1 = 0; p6_1 = 1; p7_1 = 1;
    #1 p4_1 = 0; p5_1 = 1; p6_1 = 0; p7_1 = 0;
    #1 p4_1 = 0; p5_1 = 1; p6_1 = 0; p7_1 = 1;
    #1 p4_1 = 0; p5_1 = 1; p6_1 = 1; p7_1 = 0;
    #1 p4_1 = 0; p5_1 = 1; p6_1 = 1; p7_1 = 1;
	#1 p4_1 = 1; p5_1 = 0; p6_1 = 0; p7_1 = 0;
    #1 p4_1 = 1; p5_1 = 0; p6_1 = 0; p7_1 = 1;
    #1 p4_1 = 1; p5_1 = 0; p6_1 = 1; p7_1 = 0;
    #1 p4_1 = 1; p5_1 = 0; p6_1 = 1; p7_1 = 1;
    #1 p4_1 = 1; p5_1 = 1; p6_1 = 0; p7_1 = 0;
    #1 p4_1 = 1; p5_1 = 1; p6_1 = 0; p7_1 = 1;
    #1 p4_1 = 1; p5_1 = 1; p6_1 = 1; p7_1 = 0;
    #1 p4_1 = 1; p5_1 = 1; p6_1 = 1; p7_1 = 1;
	#1 $display("");
	
  end
  
  initial begin
    #60
	$display("EJERCICIO 1: TABLA 4");
    $display("A B C D | Y");
    $display("--------|--");
    $monitor("%b %b %b %b | %b", p4_2, p5_2, p6_2, p7_2, led2_2);
       p4_2 = 0; p5_2 = 0; p6_2 = 0; p7_2 = 0;
    #1 p4_2 = 0; p5_2 = 0; p6_2 = 0; p7_2 = 1;
    #1 p4_2 = 0; p5_2 = 0; p6_2 = 1; p7_2 = 0;
    #1 p4_2 = 0; p5_2 = 0; p6_2 = 1; p7_2 = 1;
    #1 p4_2 = 0; p5_2 = 1; p6_2 = 0; p7_2 = 0;
    #1 p4_2 = 0; p5_2 = 1; p6_2 = 0; p7_2 = 1;
    #1 p4_2 = 0; p5_2 = 1; p6_2 = 1; p7_2 = 0;
    #1 p4_2 = 0; p5_2 = 1; p6_2 = 1; p7_2 = 1;
	#1 p4_2 = 1; p5_2 = 0; p6_2 = 0; p7_2 = 0;
    #1 p4_2 = 1; p5_2 = 0; p6_2 = 0; p7_2 = 1;
    #1 p4_2 = 1; p5_2 = 0; p6_2 = 1; p7_2 = 0;
    #1 p4_2 = 1; p5_2 = 0; p6_2 = 1; p7_2 = 1;
    #1 p4_2 = 1; p5_2 = 1; p6_2 = 0; p7_2 = 0;
    #1 p4_2 = 1; p5_2 = 1; p6_2 = 0; p7_2 = 1;
    #1 p4_2 = 1; p5_2 = 1; p6_2 = 1; p7_2 = 0;
    #1 p4_2 = 1; p5_2 = 1; p6_2 = 1; p7_2 = 1;
	#1 $display("");
	
  end
  
  initial begin
    #80
	$display("EJERCICIO 2: TABLA 1");
    $display("A B C D | Y");
    $display("--------|--");
    $monitor("%b %b %b %b | %b", p4_3, p5_3, p6_3, p7_3, led2_3);
       p4_3 = 0; p5_3 = 0; p6_3 = 0; p7_3 = 0;
    #1 p4_3 = 0; p5_3 = 0; p6_3 = 0; p7_3 = 1;
    #1 p4_3 = 0; p5_3 = 0; p6_3 = 1; p7_3 = 0;
    #1 p4_3 = 0; p5_3 = 0; p6_3 = 1; p7_3 = 1;
    #1 p4_3 = 0; p5_3 = 1; p6_3 = 0; p7_3 = 0;
    #1 p4_3 = 0; p5_3 = 1; p6_3 = 0; p7_3 = 1;
    #1 p4_3 = 0; p5_3 = 1; p6_3 = 1; p7_3 = 0;
    #1 p4_3 = 0; p5_3 = 1; p6_3 = 1; p7_3 = 1;
	#1 p4_3 = 1; p5_3 = 0; p6_3 = 0; p7_3 = 0;
    #1 p4_3 = 1; p5_3 = 0; p6_3 = 0; p7_3 = 1;
    #1 p4_3 = 1; p5_3 = 0; p6_3 = 1; p7_3 = 0;
    #1 p4_3 = 1; p5_3 = 0; p6_3 = 1; p7_3 = 1;
    #1 p4_3 = 1; p5_3 = 1; p6_3 = 0; p7_3 = 0;
    #1 p4_3 = 1; p5_3 = 1; p6_3 = 0; p7_3 = 1;
    #1 p4_3 = 1; p5_3 = 1; p6_3 = 1; p7_3 = 0;
    #1 p4_3 = 1; p5_3 = 1; p6_3 = 1; p7_3 = 1;
	#1 $display("");
	
  end
  
  initial begin
    #100
	$display("EJERCICIO 2: TABLA 3");
    $display("A B C D | Y");
    $display("--------|--");
    $monitor("%b %b %b %b | %b", p4_4, p5_4, p6_4, p7_4, led2_4);
       p4_4 = 0; p5_4 = 0; p6_4 = 0; p7_4 = 0;
    #1 p4_4 = 0; p5_4 = 0; p6_4 = 0; p7_4 = 1;
    #1 p4_4 = 0; p5_4 = 0; p6_4 = 1; p7_4 = 0;
    #1 p4_4 = 0; p5_4 = 0; p6_4 = 1; p7_4 = 1;
    #1 p4_4 = 0; p5_4 = 1; p6_4 = 0; p7_4 = 0;
    #1 p4_4 = 0; p5_4 = 1; p6_4 = 0; p7_4 = 1;
    #1 p4_4 = 0; p5_4 = 1; p6_4 = 1; p7_4 = 0;
    #1 p4_4 = 0; p5_4 = 1; p6_4 = 1; p7_4 = 1;
	#1 p4_4 = 1; p5_4 = 0; p6_4 = 0; p7_4 = 0;
    #1 p4_4 = 1; p5_4 = 0; p6_4 = 0; p7_4 = 1;
    #1 p4_4 = 1; p5_4 = 0; p6_4 = 1; p7_4 = 0;
    #1 p4_4 = 1; p5_4 = 0; p6_4 = 1; p7_4 = 1;
    #1 p4_4 = 1; p5_4 = 1; p6_4 = 0; p7_4 = 0;
    #1 p4_4 = 1; p5_4 = 1; p6_4 = 0; p7_4 = 1;
    #1 p4_4 = 1; p5_4 = 1; p6_4 = 1; p7_4 = 0;
    #1 p4_4 = 1; p5_4 = 1; p6_4 = 1; p7_4 = 1;
	#1 $display("");

  end
  
  initial
    #120	$finish;
  
  initial begin
    $dumpfile("Ejerccio4_tb.vcd");
    $dumpvars(0, testbench);
  end
  
endmodule